//Definicion del modulo y susu I/0
//dentro del parentesis se define los I/O

module _and(input a, input b, output c);
//2.definicion o compuertas internas
//NA
//3.Asignaciones, Intancias, Conexiones

assign C = a & b;
endmodule